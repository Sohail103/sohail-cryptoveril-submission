module stage1(
    input wire clk1,
    input wire [4:0] key_bits,
    input wire [15:0] input_data,
    output wire [15:0] stg1_out
);
    
    