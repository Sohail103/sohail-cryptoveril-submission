module stage1(key, inp, );
    